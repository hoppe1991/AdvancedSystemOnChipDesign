--------------------------------------------------------------------------------
-- filename : mips_arc_task5_btb.vhd
-- author   : Meyer zum Felde, P�ttjer, Hoppe
-- company  : TUHH
-- revision : 0.1
-- date     : 24/01/17
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

use work.mips_pkg.all;
use work.casts.all;
use work.global_pkg.all;

--------------------------------------------------------------------------------
-- Architecture of MIPS defines the pipelined MIPS (see task sheet 3) with
-- instruction cache (see task sheet 4) and BTB (see task sheet 5).
--------------------------------------------------------------------------------
architecture mips_arc_task5_btb of mips is

	-- TODO

begin
	
	-- TODO

end mips_arc_task5_btb;